library verilog;
use verilog.vl_types.all;
entity MSEND_BYTE_tb is
end MSEND_BYTE_tb;
